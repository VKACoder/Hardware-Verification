//To be updated
