//Testbench
